* Half-SRAM Core

* Library
.include "../2um_CMOS.modlib"

* MOS  D     G    S     B    MODEL  L         W
M1     nQ    BL   Vss   Vss  N_2u   l={M1_L}  w={M1_L*M1_WL}
M2     nQ    BL   Vdd   Vdd  P_2u   l={M2_L}  w={M2_L*M2_WL}
M5     nQ    WL   nBL   nBL  N_2u   l={M5_L}  w={M5_L*M5_WL}

* Cap  n1    n2   cap   ic    Rser  Lser  Cpar  m  RLShunt  temp
C1     nBL   Vss  100f

.param M1_L 2u
.param M2_L 2u
.param M5_L 2u

* Static Voltages
V1      Vdd  0   5
V5      Vss  0   0

***********************************
* Analysis 1: Finding inverter threshold
* M5 is off, so nBL can't affect this result.
* Volt  n+   n-  PULSE(V1  V2  Tdelay  Trise  Tfall  Ton  Tperiod  Ncycles)
VWL     WL   0   0
VQ      Q    0   5
VnBL    nBL  0   2.5
VBL     BL   0   0


.param M1_WL 1
.param M2_WL 3.7
.param M5_WL 1


* Estado / Precarga
.ic V(C1)=5

*.save V(nQ) V(BL) V(nBL) V(WL) V(C1)
*.step PARAM TON LIST 1.1n 1.2n 1.3n
.tran 200n


*.step param
*.step  PARAM  M2_WL LIST 1 1.5 2 2.5 3.7 5.0
*dc  Src   Vinit  Vstop  Vinc [ Src  Vinit  Vstop  Vinc ]
*.dc  VnBL  0      5      0.05

.backanno
.end
